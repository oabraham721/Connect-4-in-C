module  
    module hello_world ;
 
 initial begin
  $display ("Hello World by Deepak");
    #10  $finish;
 end

 15 endmodule // End of Module hello_world